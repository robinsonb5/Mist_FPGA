library ieee;
use ieee.numeric_std.all;

package Board_Limits is
	constant BOARD_MAX_SPRITES : integer := 52;
end package;
