//
// scandoubler_rotate.v
// 
// Copyright (c) 2024 Alastair M. Robinson
// 
// This source file is free software: you can redistribute it and/or modify 
// it under the terms of the GNU General Public License as published 
// by the Free Software Foundation, either version 3 of the License, or 
// (at your option) any later version. 
// 
// This source file is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the 
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License 
// along with this program.  If not, see <http://www.gnu.org/licenses/>. 

// Streams incoming video data to an SDRAM port, in 16-word bursts.
// Incoming data is scaled to RGB565
//
// Streams data from SDRAM to output linebuffers in 8-word bursts
// Outgoing data is scaled to OUT_COLOR_DEPTH
//
// The SDRAM controller is responsible for the actual cornerturn.
//

module scandoubler_rotate
(
	// system interface
	input        clk_sys,

	input        bypass,
	input [1:0]  rotation, // 0 - no rotation, 1 - clockwise, 2 - anticlockwise
	input        hfilter,
	input        vfilter,

	// Pixelclock
	input            pe_in,
	input            pe_out,
	input            ppe_out,

	// incoming video interface
	input        hb_in,
	input        vb_in,
	input        hs_in,
	input        vs_in,
	input [COLOR_DEPTH-1:0] r_in,
	input [COLOR_DEPTH-1:0] g_in,
	input [COLOR_DEPTH-1:0] b_in,

	// output interface
	input        hb_sd,
	input        vb_sd,
	input        vs_sd,
	output [OUT_COLOR_DEPTH-1:0] r_out,
	output [OUT_COLOR_DEPTH-1:0] g_out,
	output [OUT_COLOR_DEPTH-1:0] b_out,

	// Memory interface - to RAM.  Operates on 16-word bursts
	output reg          vidin_req,    // High at start of row, remains high until burst of 16 pixels has been delivered
	output wire         vidin_frame,  // Odd or even frame for double-buffering
	output reg [9:0]    vidin_row,    // Y position of current row.
	output reg [9:0]    vidin_col,    // X position of current burst.
	output reg [15:0]   vidin_d,      // Incoming video data
	input wire          vidin_ack,    // Request next word from host
	
	// Memory interface - from RAM.  Operates on 8-word bursts
	output wire         vidout_req,   // High at start of row, remains high until entire row has been delivered
	output wire         vidout_frame, // Odd or even frame for double-buffering
	output wire [9:0]   vidout_row,   // Y position of current row.  (Controller maintains X counter)
	output wire [9:0]   vidout_col,   // Y position of current row.  (Controller maintains X counter)
	input wire [15:0]   vidout_d,     // Outgoing video data
	input wire          vidout_ack    // Valid data available.
);

parameter HCNT_WIDTH = 10; // Resolution of scandoubler buffer
parameter COLOR_DEPTH = 6; // Bits per colour to be stored in the buffer
parameter OUT_COLOR_DEPTH = 6; // Bits per color outputted


// Scale incoming video signal to RGB565
wire [15:0] vin_rgb565;

scandoubler_scaledepth #(.IN_DEPTH(COLOR_DEPTH),.OUT_DEPTH(5)) scalein_r (.d(r_in),.q(vin_rgb565[15:11]));
scandoubler_scaledepth #(.IN_DEPTH(COLOR_DEPTH),.OUT_DEPTH(6)) scalein_g (.d(g_in),.q(vin_rgb565[10:5]));
scandoubler_scaledepth #(.IN_DEPTH(COLOR_DEPTH),.OUT_DEPTH(5)) scalein_b (.d(b_in),.q(vin_rgb565[4:0]));


// Stream incoming pixels to SDRAM, taking care of inverting either X or Y coordinates.
// The SDRAM controller does the actual cornerturn.

// Framing
reg [HCNT_WIDTH-1:0] in_xpos;
reg [HCNT_WIDTH-1:0] in_ypos=239;
reg [HCNT_WIDTH-1:0] in_xpos_max = 320;
reg [HCNT_WIDTH-1:0] in_ypos_max = 238;
reg hb_in_d;

// Toggle logical / physical frame every vblank
reg logicalframe = 1'b0;
reg vb_d = 1'b1;
reg vb_stb = 1'b0;
reg hb_stb = 1'b0;

always @(posedge clk_sys) begin
	vb_stb<=1'b0;

	vb_d<=vb_in;
	if(!vb_d && vb_in) begin
		vb_stb<=1'b1;
		logicalframe<=~logicalframe;
		in_ypos_max<=in_ypos-1'b1;
	end
end

always @(posedge clk_sys) begin
	hb_stb<=1'b0;

	hb_in_d<=hb_in;
	if(vb_in)
		in_ypos<=10'd0;
	else if(!hb_in_d && hb_in)	begin // Increment row on hblank
		hb_stb<=1'b1;
		in_ypos<=in_ypos+10'd1;
		in_xpos_max <= in_xpos;
	end
end

always @(posedge clk_sys) begin
	if(hb_in)
		in_xpos<=10'd0;
	else if(pe_in)
		in_xpos<=in_xpos+10'd1;	// Increment column on pixel enable
end

// Buffer incoming video data and write to SDRAM.
// (16 word bursts, striped across two banks, SDRAM controller handles the actual cornerturn)

reg [15:0] rowbuf[0:31] /* synthesis ramstyle="logic" */;
reg [4:0] rowwptr;
reg [4:0] rowrptr;
reg running=1'b0;

wire [3:0] escape,start;

always @(posedge clk_sys) begin

	// Reset on vblank
	if(vb_in) begin
		running<=1'b1; // (rotation!=2'b00 && !bypass);
		rowwptr<=5'h0;
	end

	// Don't update row during hblank (gives linebuffer time to empty)
	if(!hb_in) begin
		if(rotation[0])
			vidin_row<=in_ypos_max-in_ypos;
		else
			vidin_row<=in_ypos;
	end

	// Write incoming pixels to a line buffer
	if(running && pe_in && !vb_in && !hb_in) begin
		rowbuf[rowwptr]<=vin_rgb565;
		if((rowwptr[3:0]==4'b1111) || (hb_in & !hb_in_d)) begin
			vidin_col<=in_xpos;
			vidin_req<=1'b1;
			rowrptr<={rowwptr[4],4'b0000};
		end
		rowwptr<=rowwptr+1'b1;
	end

	// Write pixels from linebuffer to SDRAM
	vidin_d <= rowbuf[rowrptr];
	vidin_col[3:0] <= rowrptr[3:0];

	// Terminate burst after 16 pixels
	if(vidin_ack) begin
		if(rowrptr[3:0]==4'b1111)
			vidin_req<=1'b0;
		rowrptr<=rowrptr+1'b1;
	end
end

assign vidin_frame = logicalframe;


// Pixel read process - streams data from SDRAM to linebuffers.

reg [15:0] linebuffer1 [0:2**HCNT_WIDTH-1];
reg [15:0] linebuffer2 [0:2**HCNT_WIDTH-1];

reg fetch;

reg [HCNT_WIDTH-1:0] fetch_xpos;
reg [HCNT_WIDTH-1:0] sd_ypos;

reg hb_sd_d;
reg vs_sd_d;

reg hb_sd_stb;
reg vs_sd_stb;


// Interpolation - first calculate appropriate step size:

localparam int_fracwidth=16;
wire [HCNT_WIDTH+int_fracwidth-1:0] int_stepsize;
wire int_divdone;

unsigned_division #(.widthlog2(HCNT_WIDTH+int_fracwidth)) div (
	.clk(clk_sys),
	.reset_n(1'b1),
	.dividend({in_ypos_max[HCNT_WIDTH-2:0],{int_fracwidth+1{1'b0}}}),
	.divisor({{int_fracwidth{1'b0}},in_xpos_max}),
	.quotient(int_stepsize),
	.remainder(),
	.req(vs_sd_stb),
	.ack(int_divdone)
);

// Vertical interpolation

wire [HCNT_WIDTH-1:0] vi_whole; // Row number
wire [int_fracwidth-1:0] vi_fraction; // Blend factor
wire vi_step; // Move onto the next line
wire vi_ready;
wire vi_blank;

frac_interp #(.bitwidth(HCNT_WIDTH),.fracwidth(int_fracwidth)) interp_core_v (
	.clk(clk_sys),
	.reset_n(1'b1),
	.stepsize(int_stepsize),
	.offset(0),
	.limit(in_xpos_max),
	.step_reset(vs_sd_stb),
	.step_in(hb_sd_stb),
	.step_out(vi_step),
	.whole(vi_whole),
	.fraction(vi_fraction),
	.blank(vi_blank)
);

reg fetchbuffer;

always @(posedge clk_sys) begin
	hb_sd_stb<=1'b0;
	vs_sd_stb<=1'b0;
	hb_sd_d<=hb_sd;
	vs_sd_d<=vs_sd;

	sd_ypos <= rotation[0] ? vi_whole : in_xpos_max-vi_whole;
	
	if(!vb_sd && !hb_sd_d && hb_sd) begin // Increment row on hblank
		hb_sd_stb<=1'b1;
	end

	if (vi_step) begin
		fetch_xpos <= 10'b0;
		fetch<=1'b1;
		fetchbuffer<=fetchbuffer ^ vfilter;
	end

	if(!vs_sd_d && vs_sd) begin
		vs_sd_stb<=1'b1;
		fetch_xpos <= 10'b0;	// Pre-fetch the first row.
		fetch<=1'b1;
		fetchbuffer<=1'b0;
	end

	if(fetch && fetch_xpos==in_ypos_max)
		fetch<=1'b0;
	
	if(vidout_ack) begin
		fetch_xpos<=fetch_xpos+10'd1;
		if(fetchbuffer)
			linebuffer1[fetch_xpos]<=vidout_d;
		else
			linebuffer2[fetch_xpos]<=vidout_d;
	end
	
end

assign vidout_row = sd_ypos;
assign vidout_col = fetch_xpos;

assign vidout_frame = ~logicalframe;
assign vidout_req = fetch;


// Basic horizontal interpolation


// Offset for centering the image would be (xmax-ymax)/2
// but scandoubled high-res pixels have four times the pixel clock of original
// low-res pixels, so we use (xmax-ymax)*2.

reg [HCNT_WIDTH-1:0] hi_offset;
always @(posedge clk_sys) begin
	hi_offset<={in_xpos_max[HCNT_WIDTH-2:0],1'b0}-{in_ypos_max[HCNT_WIDTH-2:0],1'b0};
end

wire [HCNT_WIDTH-1:0] hi_whole; // Index into pixel buffer
wire [int_fracwidth-1:0] hi_fraction; // Blend factor
wire hi_step; // Move onto the next pixel
wire hi_blank;

frac_interp #(.bitwidth(HCNT_WIDTH),.fracwidth(int_fracwidth)) interp_core_h (
	.clk(clk_sys),
	.reset_n(1'b1),
	.stepsize(int_stepsize),
	.offset(hi_offset),
	.limit(in_ypos_max),
	.step_reset(hb_sd_stb),
	.step_in(!hb_sd && ppe_out),
	.step_out(hi_step),
	.whole(hi_whole),
	.fraction(hi_fraction),
	.blank(hi_blank)
);


// Interpolate pixels 

reg [7:0] hfilter_fraction;
wire [7:0] vfilter_fraction = vfilter ? vi_fraction[15:8] : 8'h00;

reg [15:0] row1_pix1;
reg [15:0] row2_pix1;
wire [15:0] col_pix1;
reg [15:0] col_pix2;
wire [15:0] final_rgb565;

reg [2:0] hi_blank_d;
reg hi_step_d;

always @(posedge clk_sys) begin
	hi_step_d<= hi_step;

	if(fetchbuffer) begin
		row1_pix1<=linebuffer1[hi_whole];
		row2_pix1<=linebuffer2[hi_whole];
	end else begin
		row2_pix1<=linebuffer1[hi_whole];
		row1_pix1<=linebuffer2[hi_whole];
	end

	// Moved this to a clock edge to keep the fraction in sync with the pixels.
	hfilter_fraction <= hfilter ? hi_fraction[15:8] : 8'h00;

	if(ppe_out)
		hi_blank_d<= {hi_blank_d[1:0],hi_blank};

	if(hi_step_d) begin
		col_pix2<=col_pix1;
	end
end

scandoubler_rgb_interp rgbinterp_v
(
	.clk_sys(clk_sys),
	.blank(vi_blank),
	.fraction(vfilter_fraction),
	.rgb_in(row1_pix1),
	.rgb_in_prev(row2_pix1),
	.rgb_out(col_pix1)
);


scandoubler_rgb_interp rgbinterp_h
(
	.clk_sys(clk_sys),
	.blank(hi_blank_d[2]),
	.fraction(hfilter_fraction),
	.rgb_in(col_pix1),
	.rgb_in_prev(col_pix2),
	.rgb_out(final_rgb565)
);

scandoubler_scaledepth #(.IN_DEPTH(5),.OUT_DEPTH(OUT_COLOR_DEPTH)) scaleout_r (.d(final_rgb565[15:11]),.q(r_out));
scandoubler_scaledepth #(.IN_DEPTH(6),.OUT_DEPTH(OUT_COLOR_DEPTH)) scaleout_g (.d(final_rgb565[10:5]),.q(g_out));
scandoubler_scaledepth #(.IN_DEPTH(5),.OUT_DEPTH(OUT_COLOR_DEPTH)) scaleout_b (.d(final_rgb565[4:0]),.q(b_out));

endmodule


